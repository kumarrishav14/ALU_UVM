`include "uvm_macros.svh"
`include "transaction.sv"
`include "dir_sequence.sv"
`include "rnd_sequence.sv"
`include "interface.sv"
`include "driver.sv"
`include "monitor.sv"
`include "agent.sv"
`include "reference_model.sv"
`include "scoreboard.sv"
`include "fun_cov.sv"
`include "environmnet.sv"
`include "test.sv"
`include "tb_top.sv"