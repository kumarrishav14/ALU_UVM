`include "uvm_macros.svh"
`include "transaction.sv"
`include "dir_sequence.sv"
`include "rnd_sequence.sv"
`include "interface.sv"
`include "driver.sv"
`include "agent.sv"
